-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb1",
     9 => x"f4080b0b",
    10 => x"0bb1f808",
    11 => x"0b0b0bb1",
    12 => x"fc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b1fc0c0b",
    16 => x"0b0bb1f8",
    17 => x"0c0b0b0b",
    18 => x"b1f40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba6f8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b1f470bc",
    57 => x"98278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"88e20402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b2840c9f",
    65 => x"0bb2880c",
    66 => x"a0717081",
    67 => x"055334b2",
    68 => x"8808ff05",
    69 => x"b2880cb2",
    70 => x"88088025",
    71 => x"eb38b284",
    72 => x"08ff05b2",
    73 => x"840cb284",
    74 => x"088025d7",
    75 => x"38800bb2",
    76 => x"880c800b",
    77 => x"b2840c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"b2840825",
    97 => x"8f3882bc",
    98 => x"2db28408",
    99 => x"ff05b284",
   100 => x"0c82fe04",
   101 => x"b28408b2",
   102 => x"88085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038b2",
   107 => x"8408a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34b28808",
   111 => x"8105b288",
   112 => x"0cb28808",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"b2880cb2",
   116 => x"84088105",
   117 => x"b2840c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134b288",
   122 => x"088105b2",
   123 => x"880cb288",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800bb288",
   127 => x"0cb28408",
   128 => x"8105b284",
   129 => x"0c028c05",
   130 => x"0d0402e8",
   131 => x"050d7779",
   132 => x"5656880b",
   133 => x"fc167771",
   134 => x"2c8f0654",
   135 => x"52548053",
   136 => x"72722595",
   137 => x"387153fb",
   138 => x"e0145187",
   139 => x"71348114",
   140 => x"ff145454",
   141 => x"72f13871",
   142 => x"53f91576",
   143 => x"712c8706",
   144 => x"53517180",
   145 => x"2e8b38fb",
   146 => x"e0145171",
   147 => x"71348114",
   148 => x"54728e24",
   149 => x"95388f73",
   150 => x"3153fbe0",
   151 => x"1451a071",
   152 => x"348114ff",
   153 => x"14545472",
   154 => x"f1380298",
   155 => x"050d0402",
   156 => x"ec050d80",
   157 => x"0bb28c0c",
   158 => x"f68c08f6",
   159 => x"90087188",
   160 => x"2c565481",
   161 => x"ff065273",
   162 => x"72258838",
   163 => x"7154820b",
   164 => x"b28c0c72",
   165 => x"882c7381",
   166 => x"ff065455",
   167 => x"7473258b",
   168 => x"3872b28c",
   169 => x"088407b2",
   170 => x"8c0c5573",
   171 => x"842b86a0",
   172 => x"71258371",
   173 => x"31700b0b",
   174 => x"0bacfc0c",
   175 => x"81712bff",
   176 => x"05f6880c",
   177 => x"fdfc13ff",
   178 => x"122c7888",
   179 => x"29ff9405",
   180 => x"70812cb2",
   181 => x"8c085258",
   182 => x"52555152",
   183 => x"5476802e",
   184 => x"85387081",
   185 => x"075170f6",
   186 => x"940c7109",
   187 => x"8105f680",
   188 => x"0c720981",
   189 => x"05f6840c",
   190 => x"0294050d",
   191 => x"0402f405",
   192 => x"0d745372",
   193 => x"70810554",
   194 => x"80f52d52",
   195 => x"71802e89",
   196 => x"38715182",
   197 => x"f82d8683",
   198 => x"04810bb1",
   199 => x"f40c028c",
   200 => x"050d0402",
   201 => x"fc050d81",
   202 => x"808051c0",
   203 => x"115170fb",
   204 => x"38028405",
   205 => x"0d0402fc",
   206 => x"050d84bf",
   207 => x"5186a32d",
   208 => x"ff115170",
   209 => x"8025f638",
   210 => x"0284050d",
   211 => x"0402fc05",
   212 => x"0dec5183",
   213 => x"710c86a3",
   214 => x"2d82710c",
   215 => x"0284050d",
   216 => x"0402fc05",
   217 => x"0dec5192",
   218 => x"710c86a3",
   219 => x"2d82710c",
   220 => x"0284050d",
   221 => x"0402d005",
   222 => x"0d7d5480",
   223 => x"5ba40bec",
   224 => x"0c7352b2",
   225 => x"90519eb6",
   226 => x"2db1f408",
   227 => x"7b2e81ab",
   228 => x"38b29408",
   229 => x"70f80c89",
   230 => x"1580f52d",
   231 => x"8a1680f5",
   232 => x"2d718280",
   233 => x"29058817",
   234 => x"80f52d70",
   235 => x"84808029",
   236 => x"12f40c7e",
   237 => x"ff155c5e",
   238 => x"57555658",
   239 => x"767b2e8b",
   240 => x"38811a77",
   241 => x"812a585a",
   242 => x"76f738f7",
   243 => x"1a5a815b",
   244 => x"80782580",
   245 => x"e6387952",
   246 => x"7651848a",
   247 => x"2db2dc52",
   248 => x"b29051a0",
   249 => x"ec2db1f4",
   250 => x"08802eb8",
   251 => x"38b2dc5c",
   252 => x"83fc597b",
   253 => x"7084055d",
   254 => x"087081ff",
   255 => x"0671882a",
   256 => x"7081ff06",
   257 => x"73902a70",
   258 => x"81ff0675",
   259 => x"982ae80c",
   260 => x"e80c58e8",
   261 => x"0c57e80c",
   262 => x"fc1a5a53",
   263 => x"788025d3",
   264 => x"3888ab04",
   265 => x"b1f4085b",
   266 => x"848058b2",
   267 => x"9051a0bf",
   268 => x"2dfc8018",
   269 => x"81185858",
   270 => x"87d00486",
   271 => x"b62d840b",
   272 => x"ec0c7a80",
   273 => x"2e8d38ad",
   274 => x"80519099",
   275 => x"2d8e9c2d",
   276 => x"88d904af",
   277 => x"c4519099",
   278 => x"2d7ab1f4",
   279 => x"0c02b005",
   280 => x"0d0402ec",
   281 => x"050d840b",
   282 => x"ec0c8dfd",
   283 => x"2d8ae72d",
   284 => x"81f72d86",
   285 => x"f551a6f3",
   286 => x"2dad8051",
   287 => x"90992d8e",
   288 => x"9c2d8af3",
   289 => x"2d90a92d",
   290 => x"ad940b80",
   291 => x"f52d7086",
   292 => x"2b80c006",
   293 => x"ada00b80",
   294 => x"f52d7087",
   295 => x"2b818006",
   296 => x"adac0b80",
   297 => x"f52d7085",
   298 => x"2ba00674",
   299 => x"730707ad",
   300 => x"b80b80f5",
   301 => x"2d708c2b",
   302 => x"80e08006",
   303 => x"adc40b80",
   304 => x"f52d7084",
   305 => x"2b900674",
   306 => x"730707ad",
   307 => x"d00b80f5",
   308 => x"2d70912b",
   309 => x"98808006",
   310 => x"addc0b80",
   311 => x"f52d708a",
   312 => x"2b988006",
   313 => x"74730707",
   314 => x"ade80b80",
   315 => x"f52d7090",
   316 => x"2b848080",
   317 => x"06adf40b",
   318 => x"80f52d70",
   319 => x"8e2b8380",
   320 => x"80067473",
   321 => x"0707ae80",
   322 => x"0b80f52d",
   323 => x"70932ba0",
   324 => x"808006ae",
   325 => x"8c0b80f5",
   326 => x"2d70942b",
   327 => x"90800a06",
   328 => x"74730707",
   329 => x"ae980b80",
   330 => x"f52d7088",
   331 => x"2b868006",
   332 => x"7207fc0c",
   333 => x"53545454",
   334 => x"54545454",
   335 => x"54545454",
   336 => x"54545454",
   337 => x"56545257",
   338 => x"57535386",
   339 => x"52b1f408",
   340 => x"8538b1f4",
   341 => x"085271ec",
   342 => x"0c898204",
   343 => x"71980c04",
   344 => x"ffb008b1",
   345 => x"f40c0481",
   346 => x"0bffb00c",
   347 => x"04800bff",
   348 => x"b00c0402",
   349 => x"f4050d8b",
   350 => x"f504b1f4",
   351 => x"0881f02e",
   352 => x"09810689",
   353 => x"38810bb0",
   354 => x"a80c8bf5",
   355 => x"04b1f408",
   356 => x"81e02e09",
   357 => x"81068938",
   358 => x"810bb0ac",
   359 => x"0c8bf504",
   360 => x"b1f40852",
   361 => x"b0ac0880",
   362 => x"2e8838b1",
   363 => x"f4088180",
   364 => x"05527184",
   365 => x"2c728f06",
   366 => x"5353b0a8",
   367 => x"08802e99",
   368 => x"38728429",
   369 => x"afe80572",
   370 => x"1381712b",
   371 => x"70097308",
   372 => x"06730c51",
   373 => x"53538beb",
   374 => x"04728429",
   375 => x"afe80572",
   376 => x"1383712b",
   377 => x"72080772",
   378 => x"0c535380",
   379 => x"0bb0ac0c",
   380 => x"800bb0a8",
   381 => x"0cb29c51",
   382 => x"8cf62db1",
   383 => x"f408ff24",
   384 => x"fef83880",
   385 => x"0bb1f40c",
   386 => x"028c050d",
   387 => x"0402f805",
   388 => x"0dafe852",
   389 => x"8f518072",
   390 => x"70840554",
   391 => x"0cff1151",
   392 => x"708025f2",
   393 => x"38028805",
   394 => x"0d0402f0",
   395 => x"050d7551",
   396 => x"8aed2d70",
   397 => x"822cfc06",
   398 => x"afe81172",
   399 => x"109e0671",
   400 => x"0870722a",
   401 => x"70830682",
   402 => x"742b7009",
   403 => x"7406760c",
   404 => x"54515657",
   405 => x"5351538a",
   406 => x"e72d71b1",
   407 => x"f40c0290",
   408 => x"050d0402",
   409 => x"fc050d72",
   410 => x"5180710c",
   411 => x"800b8412",
   412 => x"0c028405",
   413 => x"0d0402f0",
   414 => x"050d7570",
   415 => x"08841208",
   416 => x"535353ff",
   417 => x"5471712e",
   418 => x"a8388aed",
   419 => x"2d841308",
   420 => x"70842914",
   421 => x"88117008",
   422 => x"7081ff06",
   423 => x"84180881",
   424 => x"11870684",
   425 => x"1a0c5351",
   426 => x"55515151",
   427 => x"8ae72d71",
   428 => x"5473b1f4",
   429 => x"0c029005",
   430 => x"0d0402f8",
   431 => x"050d8aed",
   432 => x"2de00870",
   433 => x"8b2a7081",
   434 => x"06515252",
   435 => x"70802e9d",
   436 => x"38b29c08",
   437 => x"708429b2",
   438 => x"a4057381",
   439 => x"ff06710c",
   440 => x"5151b29c",
   441 => x"08811187",
   442 => x"06b29c0c",
   443 => x"51800bb2",
   444 => x"c40c8ae0",
   445 => x"2d8ae72d",
   446 => x"0288050d",
   447 => x"0402fc05",
   448 => x"0db29c51",
   449 => x"8ce32d8c",
   450 => x"8d2d8dba",
   451 => x"518adc2d",
   452 => x"0284050d",
   453 => x"04b2c808",
   454 => x"b1f40c04",
   455 => x"02fc050d",
   456 => x"8ea6048a",
   457 => x"f32d80f6",
   458 => x"518caa2d",
   459 => x"b1f408f3",
   460 => x"3880da51",
   461 => x"8caa2db1",
   462 => x"f408e838",
   463 => x"b1f408b0",
   464 => x"b40cb1f4",
   465 => x"085184ef",
   466 => x"2d028405",
   467 => x"0d0402ec",
   468 => x"050d7654",
   469 => x"8052870b",
   470 => x"881580f5",
   471 => x"2d565374",
   472 => x"72248338",
   473 => x"a0537251",
   474 => x"82f82d81",
   475 => x"128b1580",
   476 => x"f52d5452",
   477 => x"727225de",
   478 => x"38029405",
   479 => x"0d0402f0",
   480 => x"050db2c8",
   481 => x"085481f7",
   482 => x"2d800bb2",
   483 => x"cc0c7308",
   484 => x"802e8180",
   485 => x"38820bb2",
   486 => x"880cb2cc",
   487 => x"088f06b2",
   488 => x"840c7308",
   489 => x"5271832e",
   490 => x"96387183",
   491 => x"26893871",
   492 => x"812eaf38",
   493 => x"8fff0471",
   494 => x"852e9f38",
   495 => x"8fff0488",
   496 => x"1480f52d",
   497 => x"841508ac",
   498 => x"94535452",
   499 => x"85fd2d71",
   500 => x"84291370",
   501 => x"08525290",
   502 => x"83047351",
   503 => x"8ece2d8f",
   504 => x"ff04b0b0",
   505 => x"08881508",
   506 => x"2c708106",
   507 => x"51527180",
   508 => x"2e8738ac",
   509 => x"98518ffc",
   510 => x"04ac9c51",
   511 => x"85fd2d84",
   512 => x"14085185",
   513 => x"fd2db2cc",
   514 => x"088105b2",
   515 => x"cc0c8c14",
   516 => x"548f8e04",
   517 => x"0290050d",
   518 => x"0471b2c8",
   519 => x"0c8efe2d",
   520 => x"b2cc08ff",
   521 => x"05b2d00c",
   522 => x"0402e805",
   523 => x"0db2c808",
   524 => x"b2d40857",
   525 => x"5587518c",
   526 => x"aa2db1f4",
   527 => x"08812a70",
   528 => x"81065152",
   529 => x"71802ea0",
   530 => x"3890cf04",
   531 => x"8af32d87",
   532 => x"518caa2d",
   533 => x"b1f408f4",
   534 => x"38b0b408",
   535 => x"813270b0",
   536 => x"b40c7052",
   537 => x"5284ef2d",
   538 => x"80fe518c",
   539 => x"aa2db1f4",
   540 => x"08802ea6",
   541 => x"38b0b408",
   542 => x"802e9138",
   543 => x"800bb0b4",
   544 => x"0c805184",
   545 => x"ef2d918c",
   546 => x"048af32d",
   547 => x"80fe518c",
   548 => x"aa2db1f4",
   549 => x"08f33886",
   550 => x"e12db0b4",
   551 => x"08903881",
   552 => x"fd518caa",
   553 => x"2d81fa51",
   554 => x"8caa2d96",
   555 => x"df0481f5",
   556 => x"518caa2d",
   557 => x"b1f40881",
   558 => x"2a708106",
   559 => x"51527180",
   560 => x"2eaf38b2",
   561 => x"d0085271",
   562 => x"802e8938",
   563 => x"ff12b2d0",
   564 => x"0c91f104",
   565 => x"b2cc0810",
   566 => x"b2cc0805",
   567 => x"70842916",
   568 => x"51528812",
   569 => x"08802e89",
   570 => x"38ff5188",
   571 => x"12085271",
   572 => x"2d81f251",
   573 => x"8caa2db1",
   574 => x"f408812a",
   575 => x"70810651",
   576 => x"5271802e",
   577 => x"b138b2cc",
   578 => x"08ff11b2",
   579 => x"d0085653",
   580 => x"53737225",
   581 => x"89388114",
   582 => x"b2d00c92",
   583 => x"b6047210",
   584 => x"13708429",
   585 => x"16515288",
   586 => x"1208802e",
   587 => x"8938fe51",
   588 => x"88120852",
   589 => x"712d81fd",
   590 => x"518caa2d",
   591 => x"b1f40881",
   592 => x"2a708106",
   593 => x"51527180",
   594 => x"2ead38b2",
   595 => x"d008802e",
   596 => x"8938800b",
   597 => x"b2d00c92",
   598 => x"f704b2cc",
   599 => x"0810b2cc",
   600 => x"08057084",
   601 => x"29165152",
   602 => x"88120880",
   603 => x"2e8938fd",
   604 => x"51881208",
   605 => x"52712d81",
   606 => x"fa518caa",
   607 => x"2db1f408",
   608 => x"812a7081",
   609 => x"06515271",
   610 => x"802eae38",
   611 => x"b2cc08ff",
   612 => x"115452b2",
   613 => x"d0087325",
   614 => x"883872b2",
   615 => x"d00c93b9",
   616 => x"04711012",
   617 => x"70842916",
   618 => x"51528812",
   619 => x"08802e89",
   620 => x"38fc5188",
   621 => x"12085271",
   622 => x"2db2d008",
   623 => x"70535473",
   624 => x"802e8a38",
   625 => x"8c15ff15",
   626 => x"555593bf",
   627 => x"04820bb2",
   628 => x"880c718f",
   629 => x"06b2840c",
   630 => x"81eb518c",
   631 => x"aa2db1f4",
   632 => x"08812a70",
   633 => x"81065152",
   634 => x"71802ead",
   635 => x"38740885",
   636 => x"2e098106",
   637 => x"a4388815",
   638 => x"80f52dff",
   639 => x"05527188",
   640 => x"1681b72d",
   641 => x"71982b52",
   642 => x"71802588",
   643 => x"38800b88",
   644 => x"1681b72d",
   645 => x"74518ece",
   646 => x"2d81f451",
   647 => x"8caa2db1",
   648 => x"f408812a",
   649 => x"70810651",
   650 => x"5271802e",
   651 => x"b3387408",
   652 => x"852e0981",
   653 => x"06aa3888",
   654 => x"1580f52d",
   655 => x"81055271",
   656 => x"881681b7",
   657 => x"2d7181ff",
   658 => x"068b1680",
   659 => x"f52d5452",
   660 => x"72722787",
   661 => x"38728816",
   662 => x"81b72d74",
   663 => x"518ece2d",
   664 => x"80da518c",
   665 => x"aa2db1f4",
   666 => x"08812a70",
   667 => x"81065152",
   668 => x"71802e81",
   669 => x"a638b2c8",
   670 => x"08b2d008",
   671 => x"55537380",
   672 => x"2e8a388c",
   673 => x"13ff1555",
   674 => x"5394fe04",
   675 => x"72085271",
   676 => x"822ea638",
   677 => x"71822689",
   678 => x"3871812e",
   679 => x"a938969b",
   680 => x"0471832e",
   681 => x"b1387184",
   682 => x"2e098106",
   683 => x"80ed3888",
   684 => x"13085190",
   685 => x"992d969b",
   686 => x"04b2d008",
   687 => x"51881308",
   688 => x"52712d96",
   689 => x"9b04810b",
   690 => x"8814082b",
   691 => x"b0b00832",
   692 => x"b0b00c95",
   693 => x"f1048813",
   694 => x"80f52d81",
   695 => x"058b1480",
   696 => x"f52d5354",
   697 => x"71742483",
   698 => x"38805473",
   699 => x"881481b7",
   700 => x"2d8efe2d",
   701 => x"969b0475",
   702 => x"08802ea2",
   703 => x"38750851",
   704 => x"8caa2db1",
   705 => x"f4088106",
   706 => x"5271802e",
   707 => x"8b38b2d0",
   708 => x"08518416",
   709 => x"0852712d",
   710 => x"88165675",
   711 => x"da388054",
   712 => x"800bb288",
   713 => x"0c738f06",
   714 => x"b2840ca0",
   715 => x"5273b2d0",
   716 => x"082e0981",
   717 => x"069838b2",
   718 => x"cc08ff05",
   719 => x"74327009",
   720 => x"81057072",
   721 => x"079f2a91",
   722 => x"71315151",
   723 => x"53537151",
   724 => x"82f82d81",
   725 => x"14548e74",
   726 => x"25c638b0",
   727 => x"b4085271",
   728 => x"b1f40c02",
   729 => x"98050d04",
   730 => x"02f4050d",
   731 => x"d45281ff",
   732 => x"720c7108",
   733 => x"5381ff72",
   734 => x"0c72882b",
   735 => x"83fe8006",
   736 => x"72087081",
   737 => x"ff065152",
   738 => x"5381ff72",
   739 => x"0c727107",
   740 => x"882b7208",
   741 => x"7081ff06",
   742 => x"51525381",
   743 => x"ff720c72",
   744 => x"7107882b",
   745 => x"72087081",
   746 => x"ff067207",
   747 => x"b1f40c52",
   748 => x"53028c05",
   749 => x"0d0402f4",
   750 => x"050d7476",
   751 => x"7181ff06",
   752 => x"d40c5353",
   753 => x"b2d80885",
   754 => x"3871892b",
   755 => x"5271982a",
   756 => x"d40c7190",
   757 => x"2a7081ff",
   758 => x"06d40c51",
   759 => x"71882a70",
   760 => x"81ff06d4",
   761 => x"0c517181",
   762 => x"ff06d40c",
   763 => x"72902a70",
   764 => x"81ff06d4",
   765 => x"0c51d408",
   766 => x"7081ff06",
   767 => x"515182b8",
   768 => x"bf527081",
   769 => x"ff2e0981",
   770 => x"06943881",
   771 => x"ff0bd40c",
   772 => x"d4087081",
   773 => x"ff06ff14",
   774 => x"54515171",
   775 => x"e53870b1",
   776 => x"f40c028c",
   777 => x"050d0402",
   778 => x"e8050d78",
   779 => x"55805681",
   780 => x"ff0bd40c",
   781 => x"d008708f",
   782 => x"2a708106",
   783 => x"51515372",
   784 => x"f3388281",
   785 => x"0bd00c81",
   786 => x"ff0bd40c",
   787 => x"775287fc",
   788 => x"80d15197",
   789 => x"b62d80db",
   790 => x"c6df54b1",
   791 => x"f408802e",
   792 => x"8a38ace4",
   793 => x"5185fd2d",
   794 => x"99be0481",
   795 => x"ff0bd40c",
   796 => x"d4087081",
   797 => x"ff065153",
   798 => x"7281fe2e",
   799 => x"0981069d",
   800 => x"3880ff53",
   801 => x"96e82db1",
   802 => x"f4087570",
   803 => x"8405570c",
   804 => x"ff135372",
   805 => x"8025ed38",
   806 => x"815699a3",
   807 => x"04ff1454",
   808 => x"73c93881",
   809 => x"ff0bd40c",
   810 => x"81ff0bd4",
   811 => x"0cd00870",
   812 => x"8f2a7081",
   813 => x"06515153",
   814 => x"72f33872",
   815 => x"d00c75b1",
   816 => x"f40c0298",
   817 => x"050d0402",
   818 => x"e8050d77",
   819 => x"797b5855",
   820 => x"55805372",
   821 => x"7625a338",
   822 => x"74708105",
   823 => x"5680f52d",
   824 => x"74708105",
   825 => x"5680f52d",
   826 => x"52527171",
   827 => x"2e863881",
   828 => x"5199fc04",
   829 => x"81135399",
   830 => x"d3048051",
   831 => x"70b1f40c",
   832 => x"0298050d",
   833 => x"0402ec05",
   834 => x"0d765574",
   835 => x"802ebb38",
   836 => x"9a1580e0",
   837 => x"2d51a1c2",
   838 => x"2db1f408",
   839 => x"b1f408b9",
   840 => x"840cb1f4",
   841 => x"085454b8",
   842 => x"e808802e",
   843 => x"99389415",
   844 => x"80e02d51",
   845 => x"a1c22db1",
   846 => x"f408902b",
   847 => x"83fff00a",
   848 => x"06707507",
   849 => x"515372b9",
   850 => x"840cb984",
   851 => x"08537280",
   852 => x"2e9938b8",
   853 => x"e008fe14",
   854 => x"7129b8f4",
   855 => x"0805b988",
   856 => x"0c70842b",
   857 => x"b8ec0c54",
   858 => x"9b9104b8",
   859 => x"f808b984",
   860 => x"0cb8fc08",
   861 => x"b9880cb8",
   862 => x"e808802e",
   863 => x"8a38b8e0",
   864 => x"08842b53",
   865 => x"9b8d04b9",
   866 => x"8008842b",
   867 => x"5372b8ec",
   868 => x"0c029405",
   869 => x"0d0402ec",
   870 => x"050d7670",
   871 => x"872c7180",
   872 => x"ff065556",
   873 => x"54b8e808",
   874 => x"8a387388",
   875 => x"2c7481ff",
   876 => x"065455b2",
   877 => x"dc52b8f0",
   878 => x"08155198",
   879 => x"a72db1f4",
   880 => x"0854b1f4",
   881 => x"08802eb3",
   882 => x"38b8e808",
   883 => x"802e9838",
   884 => x"728429b2",
   885 => x"dc057008",
   886 => x"5253a192",
   887 => x"2db1f408",
   888 => x"f00a0653",
   889 => x"9bf90472",
   890 => x"10b2dc05",
   891 => x"7080e02d",
   892 => x"5253a1c2",
   893 => x"2db1f408",
   894 => x"53725473",
   895 => x"b1f40c02",
   896 => x"94050d04",
   897 => x"02e0050d",
   898 => x"7970842c",
   899 => x"b9880805",
   900 => x"718f0652",
   901 => x"55537289",
   902 => x"38b2dc52",
   903 => x"735198a7",
   904 => x"2d72a029",
   905 => x"b2dc0554",
   906 => x"807480f5",
   907 => x"2d565374",
   908 => x"732e8338",
   909 => x"81537481",
   910 => x"e52e81ef",
   911 => x"38817074",
   912 => x"06545872",
   913 => x"802e81e3",
   914 => x"388b1480",
   915 => x"f52d7083",
   916 => x"2a790658",
   917 => x"56769838",
   918 => x"b0b80853",
   919 => x"72883872",
   920 => x"b6dc0b81",
   921 => x"b72d76b0",
   922 => x"b80c7353",
   923 => x"9ead0475",
   924 => x"8f2e0981",
   925 => x"0681b438",
   926 => x"749f068d",
   927 => x"29b6cf11",
   928 => x"51538114",
   929 => x"80f52d73",
   930 => x"70810555",
   931 => x"81b72d83",
   932 => x"1480f52d",
   933 => x"73708105",
   934 => x"5581b72d",
   935 => x"851480f5",
   936 => x"2d737081",
   937 => x"055581b7",
   938 => x"2d871480",
   939 => x"f52d7370",
   940 => x"81055581",
   941 => x"b72d8914",
   942 => x"80f52d73",
   943 => x"70810555",
   944 => x"81b72d8e",
   945 => x"1480f52d",
   946 => x"73708105",
   947 => x"5581b72d",
   948 => x"901480f5",
   949 => x"2d737081",
   950 => x"055581b7",
   951 => x"2d921480",
   952 => x"f52d7370",
   953 => x"81055581",
   954 => x"b72d9414",
   955 => x"80f52d73",
   956 => x"70810555",
   957 => x"81b72d96",
   958 => x"1480f52d",
   959 => x"73708105",
   960 => x"5581b72d",
   961 => x"981480f5",
   962 => x"2d737081",
   963 => x"055581b7",
   964 => x"2d9c1480",
   965 => x"f52d7370",
   966 => x"81055581",
   967 => x"b72d9e14",
   968 => x"80f52d73",
   969 => x"81b72d77",
   970 => x"b0b80c80",
   971 => x"5372b1f4",
   972 => x"0c02a005",
   973 => x"0d0402cc",
   974 => x"050d7e60",
   975 => x"5e5a800b",
   976 => x"b98408b9",
   977 => x"8808595c",
   978 => x"568058b8",
   979 => x"ec08782e",
   980 => x"81ae3877",
   981 => x"8f06a017",
   982 => x"5754738f",
   983 => x"38b2dc52",
   984 => x"76518117",
   985 => x"5798a72d",
   986 => x"b2dc5680",
   987 => x"7680f52d",
   988 => x"56547474",
   989 => x"2e833881",
   990 => x"547481e5",
   991 => x"2e80f638",
   992 => x"81707506",
   993 => x"555c7380",
   994 => x"2e80ea38",
   995 => x"8b1680f5",
   996 => x"2d980659",
   997 => x"7880de38",
   998 => x"8b537c52",
   999 => x"755199c7",
  1000 => x"2db1f408",
  1001 => x"80cf389c",
  1002 => x"160851a1",
  1003 => x"922db1f4",
  1004 => x"08841b0c",
  1005 => x"9a1680e0",
  1006 => x"2d51a1c2",
  1007 => x"2db1f408",
  1008 => x"b1f40888",
  1009 => x"1c0cb1f4",
  1010 => x"085555b8",
  1011 => x"e808802e",
  1012 => x"98389416",
  1013 => x"80e02d51",
  1014 => x"a1c22db1",
  1015 => x"f408902b",
  1016 => x"83fff00a",
  1017 => x"06701651",
  1018 => x"5473881b",
  1019 => x"0c787a0c",
  1020 => x"7b54a0b6",
  1021 => x"04811858",
  1022 => x"b8ec0878",
  1023 => x"26fed438",
  1024 => x"b8e80880",
  1025 => x"2eae387a",
  1026 => x"519b962d",
  1027 => x"b1f408b1",
  1028 => x"f40880ff",
  1029 => x"fffff806",
  1030 => x"555b7380",
  1031 => x"fffffff8",
  1032 => x"2e9238b1",
  1033 => x"f408fe05",
  1034 => x"b8e00829",
  1035 => x"b8f40805",
  1036 => x"579ec904",
  1037 => x"805473b1",
  1038 => x"f40c02b4",
  1039 => x"050d0402",
  1040 => x"f4050d74",
  1041 => x"70088105",
  1042 => x"710c7008",
  1043 => x"b8e40806",
  1044 => x"5353718e",
  1045 => x"38881308",
  1046 => x"519b962d",
  1047 => x"b1f40888",
  1048 => x"140c810b",
  1049 => x"b1f40c02",
  1050 => x"8c050d04",
  1051 => x"02f0050d",
  1052 => x"75881108",
  1053 => x"fe05b8e0",
  1054 => x"0829b8f4",
  1055 => x"08117208",
  1056 => x"b8e40806",
  1057 => x"05795553",
  1058 => x"545498a7",
  1059 => x"2d029005",
  1060 => x"0d0402f4",
  1061 => x"050d7470",
  1062 => x"882a83fe",
  1063 => x"80067072",
  1064 => x"982a0772",
  1065 => x"882b87fc",
  1066 => x"80800673",
  1067 => x"982b81f0",
  1068 => x"0a067173",
  1069 => x"0707b1f4",
  1070 => x"0c565153",
  1071 => x"51028c05",
  1072 => x"0d0402f8",
  1073 => x"050d028e",
  1074 => x"0580f52d",
  1075 => x"74882b07",
  1076 => x"7083ffff",
  1077 => x"06b1f40c",
  1078 => x"51028805",
  1079 => x"0d0402f4",
  1080 => x"050d7476",
  1081 => x"78535452",
  1082 => x"80712597",
  1083 => x"38727081",
  1084 => x"055480f5",
  1085 => x"2d727081",
  1086 => x"055481b7",
  1087 => x"2dff1151",
  1088 => x"70eb3880",
  1089 => x"7281b72d",
  1090 => x"028c050d",
  1091 => x"0402e805",
  1092 => x"0d775680",
  1093 => x"70565473",
  1094 => x"7624b138",
  1095 => x"b8ec0874",
  1096 => x"2eaa3873",
  1097 => x"519c842d",
  1098 => x"b1f408b1",
  1099 => x"f4080981",
  1100 => x"0570b1f4",
  1101 => x"08079f2a",
  1102 => x"77058117",
  1103 => x"57575353",
  1104 => x"74762488",
  1105 => x"38b8ec08",
  1106 => x"7426d838",
  1107 => x"72b1f40c",
  1108 => x"0298050d",
  1109 => x"0402f005",
  1110 => x"0db1f008",
  1111 => x"1651a28d",
  1112 => x"2db1f408",
  1113 => x"802e9b38",
  1114 => x"8b53b1f4",
  1115 => x"0852b6dc",
  1116 => x"51a1de2d",
  1117 => x"b98c0854",
  1118 => x"73802e86",
  1119 => x"38b6dc51",
  1120 => x"732d0290",
  1121 => x"050d0402",
  1122 => x"dc050d80",
  1123 => x"705a5574",
  1124 => x"b1f00825",
  1125 => x"af38b8ec",
  1126 => x"08752ea8",
  1127 => x"3878519c",
  1128 => x"842db1f4",
  1129 => x"08098105",
  1130 => x"70b1f408",
  1131 => x"079f2a76",
  1132 => x"05811b5b",
  1133 => x"565474b1",
  1134 => x"f0082588",
  1135 => x"38b8ec08",
  1136 => x"7926da38",
  1137 => x"805578b8",
  1138 => x"ec082781",
  1139 => x"cd387851",
  1140 => x"9c842db1",
  1141 => x"f408802e",
  1142 => x"81a238b1",
  1143 => x"f4088b05",
  1144 => x"80f52d70",
  1145 => x"842a7081",
  1146 => x"06771078",
  1147 => x"842bb6dc",
  1148 => x"0b80f52d",
  1149 => x"5c5c5351",
  1150 => x"55567380",
  1151 => x"2e80c638",
  1152 => x"7416822b",
  1153 => x"a5bd0bb0",
  1154 => x"c4120c54",
  1155 => x"77753110",
  1156 => x"b9901155",
  1157 => x"56907470",
  1158 => x"81055681",
  1159 => x"b72da074",
  1160 => x"81b72d76",
  1161 => x"81ff0681",
  1162 => x"16585473",
  1163 => x"802e8938",
  1164 => x"9c53b6dc",
  1165 => x"52a4be04",
  1166 => x"8b53b1f4",
  1167 => x"0852b992",
  1168 => x"1651a4f4",
  1169 => x"04741682",
  1170 => x"2ba2d50b",
  1171 => x"b0c4120c",
  1172 => x"547681ff",
  1173 => x"06811658",
  1174 => x"5473802e",
  1175 => x"89389c53",
  1176 => x"b6dc52a4",
  1177 => x"ec048b53",
  1178 => x"b1f40852",
  1179 => x"77753110",
  1180 => x"b9900551",
  1181 => x"7655a1de",
  1182 => x"2da58f04",
  1183 => x"74902975",
  1184 => x"317010b9",
  1185 => x"90055154",
  1186 => x"b1f40874",
  1187 => x"81b72d81",
  1188 => x"1959748b",
  1189 => x"24a238a3",
  1190 => x"c6047490",
  1191 => x"29753170",
  1192 => x"10b99005",
  1193 => x"8c773157",
  1194 => x"51548074",
  1195 => x"81b72d9e",
  1196 => x"14ff1656",
  1197 => x"5474f338",
  1198 => x"02a4050d",
  1199 => x"0402fc05",
  1200 => x"0db1f008",
  1201 => x"1351a28d",
  1202 => x"2db1f408",
  1203 => x"802e8838",
  1204 => x"b1f40851",
  1205 => x"9a852d80",
  1206 => x"0bb1f00c",
  1207 => x"a3872d8e",
  1208 => x"fe2d0284",
  1209 => x"050d0402",
  1210 => x"fc050d72",
  1211 => x"5170fd2e",
  1212 => x"ad3870fd",
  1213 => x"248a3870",
  1214 => x"fc2e80c4",
  1215 => x"38a6c804",
  1216 => x"70fe2eb1",
  1217 => x"3870ff2e",
  1218 => x"098106bc",
  1219 => x"38b1f008",
  1220 => x"5170802e",
  1221 => x"b338ff11",
  1222 => x"b1f00ca6",
  1223 => x"c804b1f0",
  1224 => x"08f00570",
  1225 => x"b1f00c51",
  1226 => x"7080259c",
  1227 => x"38800bb1",
  1228 => x"f00ca6c8",
  1229 => x"04b1f008",
  1230 => x"8105b1f0",
  1231 => x"0ca6c804",
  1232 => x"b1f00890",
  1233 => x"05b1f00c",
  1234 => x"a3872d8e",
  1235 => x"fe2d0284",
  1236 => x"050d0402",
  1237 => x"fc050d80",
  1238 => x"0bb1f00c",
  1239 => x"a3872d8e",
  1240 => x"952db1f4",
  1241 => x"08b1e00c",
  1242 => x"b0bc5190",
  1243 => x"992d0284",
  1244 => x"050d0471",
  1245 => x"b98c0c04",
  1246 => x"00ffffff",
  1247 => x"ff00ffff",
  1248 => x"ffff00ff",
  1249 => x"ffffff00",
  1250 => x"52657365",
  1251 => x"74000000",
  1252 => x"43617267",
  1253 => x"6172204d",
  1254 => x"6564696f",
  1255 => x"20100000",
  1256 => x"45786974",
  1257 => x"00000000",
  1258 => x"4a6f7973",
  1259 => x"7469636b",
  1260 => x"20437572",
  1261 => x"736f7200",
  1262 => x"4a6f7973",
  1263 => x"7469636b",
  1264 => x"2053696e",
  1265 => x"636c6169",
  1266 => x"72000000",
  1267 => x"4a6f7973",
  1268 => x"7469636b",
  1269 => x"205a5838",
  1270 => x"31000000",
  1271 => x"4368726f",
  1272 => x"6d613831",
  1273 => x"20446573",
  1274 => x"61637469",
  1275 => x"7661646f",
  1276 => x"00000000",
  1277 => x"4368726f",
  1278 => x"6d613831",
  1279 => x"20416374",
  1280 => x"69766164",
  1281 => x"6f000000",
  1282 => x"51532043",
  1283 => x"48525320",
  1284 => x"41637469",
  1285 => x"7661646f",
  1286 => x"28463129",
  1287 => x"00000000",
  1288 => x"51532043",
  1289 => x"48525320",
  1290 => x"44657361",
  1291 => x"63746976",
  1292 => x"61646f00",
  1293 => x"43485224",
  1294 => x"3132382f",
  1295 => x"55444720",
  1296 => x"31323820",
  1297 => x"43686172",
  1298 => x"73000000",
  1299 => x"43485224",
  1300 => x"3132382f",
  1301 => x"55444720",
  1302 => x"36342043",
  1303 => x"68617273",
  1304 => x"00000000",
  1305 => x"43485224",
  1306 => x"3132382f",
  1307 => x"55444720",
  1308 => x"44657361",
  1309 => x"63746976",
  1310 => x"61646f00",
  1311 => x"52414d20",
  1312 => x"42616a61",
  1313 => x"204f6666",
  1314 => x"00000000",
  1315 => x"52414d20",
  1316 => x"42616a61",
  1317 => x"20384b42",
  1318 => x"00000000",
  1319 => x"52414d20",
  1320 => x"5072696e",
  1321 => x"63697061",
  1322 => x"6c203136",
  1323 => x"4b420000",
  1324 => x"52414d20",
  1325 => x"5072696e",
  1326 => x"63697061",
  1327 => x"6c203332",
  1328 => x"4b420000",
  1329 => x"52414d20",
  1330 => x"5072696e",
  1331 => x"63697061",
  1332 => x"6c203438",
  1333 => x"4b420000",
  1334 => x"52414d20",
  1335 => x"5072696e",
  1336 => x"63697061",
  1337 => x"6c20314b",
  1338 => x"42000000",
  1339 => x"56656c6f",
  1340 => x"63696461",
  1341 => x"64204f72",
  1342 => x"6967696e",
  1343 => x"616c0000",
  1344 => x"56656c6f",
  1345 => x"63696461",
  1346 => x"64204e6f",
  1347 => x"57616974",
  1348 => x"00000000",
  1349 => x"56656c6f",
  1350 => x"63696461",
  1351 => x"64207832",
  1352 => x"00000000",
  1353 => x"56656c6f",
  1354 => x"63696461",
  1355 => x"64207838",
  1356 => x"00000000",
  1357 => x"5a583831",
  1358 => x"00000000",
  1359 => x"5a583830",
  1360 => x"00000000",
  1361 => x"5363616e",
  1362 => x"6c696e65",
  1363 => x"73204e6f",
  1364 => x"6e650000",
  1365 => x"5363616e",
  1366 => x"6c696e65",
  1367 => x"73204352",
  1368 => x"54203235",
  1369 => x"25000000",
  1370 => x"5363616e",
  1371 => x"6c696e65",
  1372 => x"73204352",
  1373 => x"54203530",
  1374 => x"25000000",
  1375 => x"5363616e",
  1376 => x"6c696e65",
  1377 => x"73204352",
  1378 => x"54203735",
  1379 => x"25000000",
  1380 => x"426f7264",
  1381 => x"65204e65",
  1382 => x"67726f20",
  1383 => x"4f666600",
  1384 => x"426f7264",
  1385 => x"65204e65",
  1386 => x"67726f20",
  1387 => x"4f6e0000",
  1388 => x"56696465",
  1389 => x"6f20496e",
  1390 => x"7665736f",
  1391 => x"204f6666",
  1392 => x"00000000",
  1393 => x"56696465",
  1394 => x"6f20496e",
  1395 => x"7665736f",
  1396 => x"204f6e00",
  1397 => x"56696465",
  1398 => x"6f204672",
  1399 => x"65712035",
  1400 => x"30487a00",
  1401 => x"56696465",
  1402 => x"6f204672",
  1403 => x"65712036",
  1404 => x"30487a00",
  1405 => x"50656e74",
  1406 => x"61676f6e",
  1407 => x"00000000",
  1408 => x"43617267",
  1409 => x"61204661",
  1410 => x"6c6c6964",
  1411 => x"61000000",
  1412 => x"4f4b0000",
  1413 => x"16200000",
  1414 => x"14200000",
  1415 => x"15200000",
  1416 => x"53442069",
  1417 => x"6e69742e",
  1418 => x"2e2e0a00",
  1419 => x"53442063",
  1420 => x"61726420",
  1421 => x"72657365",
  1422 => x"74206661",
  1423 => x"696c6564",
  1424 => x"210a0000",
  1425 => x"53444843",
  1426 => x"20657272",
  1427 => x"6f72210a",
  1428 => x"00000000",
  1429 => x"57726974",
  1430 => x"65206661",
  1431 => x"696c6564",
  1432 => x"0a000000",
  1433 => x"52656164",
  1434 => x"20666169",
  1435 => x"6c65640a",
  1436 => x"00000000",
  1437 => x"4261636b",
  1438 => x"00000000",
  1439 => x"00000002",
  1440 => x"00000002",
  1441 => x"00001388",
  1442 => x"0000034d",
  1443 => x"00000003",
  1444 => x"000017b8",
  1445 => x"00000002",
  1446 => x"00000003",
  1447 => x"000017b0",
  1448 => x"00000002",
  1449 => x"00000003",
  1450 => x"000017a8",
  1451 => x"00000002",
  1452 => x"00000003",
  1453 => x"00001798",
  1454 => x"00000004",
  1455 => x"00000003",
  1456 => x"00001790",
  1457 => x"00000002",
  1458 => x"00000003",
  1459 => x"00001780",
  1460 => x"00000004",
  1461 => x"00000003",
  1462 => x"00001770",
  1463 => x"00000004",
  1464 => x"00000003",
  1465 => x"00001768",
  1466 => x"00000002",
  1467 => x"00000003",
  1468 => x"0000175c",
  1469 => x"00000003",
  1470 => x"00000003",
  1471 => x"00001754",
  1472 => x"00000002",
  1473 => x"00000003",
  1474 => x"0000174c",
  1475 => x"00000002",
  1476 => x"00000003",
  1477 => x"00001740",
  1478 => x"00000003",
  1479 => x"00000002",
  1480 => x"00001390",
  1481 => x"00001353",
  1482 => x"00000002",
  1483 => x"000013a0",
  1484 => x"0000071c",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"000013a8",
  1489 => x"000013b8",
  1490 => x"000013cc",
  1491 => x"000013dc",
  1492 => x"000013f4",
  1493 => x"00001408",
  1494 => x"00001420",
  1495 => x"00001434",
  1496 => x"0000144c",
  1497 => x"00001464",
  1498 => x"0000147c",
  1499 => x"0000148c",
  1500 => x"0000149c",
  1501 => x"000014b0",
  1502 => x"000014c4",
  1503 => x"000014d8",
  1504 => x"000014ec",
  1505 => x"00001500",
  1506 => x"00001514",
  1507 => x"00001524",
  1508 => x"00001534",
  1509 => x"0000153c",
  1510 => x"00001544",
  1511 => x"00001554",
  1512 => x"00001568",
  1513 => x"0000157c",
  1514 => x"00001590",
  1515 => x"000015a0",
  1516 => x"000015b0",
  1517 => x"000015c4",
  1518 => x"000015d4",
  1519 => x"000015e4",
  1520 => x"000015f4",
  1521 => x"00000004",
  1522 => x"00001600",
  1523 => x"000017c4",
  1524 => x"00000004",
  1525 => x"00001610",
  1526 => x"00001680",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000000",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
  1539 => x"00000000",
  1540 => x"00000000",
  1541 => x"00000000",
  1542 => x"00000000",
  1543 => x"00000000",
  1544 => x"00000000",
  1545 => x"00000000",
  1546 => x"00000000",
  1547 => x"00000000",
  1548 => x"00000000",
  1549 => x"00000000",
  1550 => x"00000000",
  1551 => x"00000002",
  1552 => x"00001c90",
  1553 => x"00001155",
  1554 => x"00000002",
  1555 => x"00001cae",
  1556 => x"00001155",
  1557 => x"00000002",
  1558 => x"00001ccc",
  1559 => x"00001155",
  1560 => x"00000002",
  1561 => x"00001cea",
  1562 => x"00001155",
  1563 => x"00000002",
  1564 => x"00001d08",
  1565 => x"00001155",
  1566 => x"00000002",
  1567 => x"00001d26",
  1568 => x"00001155",
  1569 => x"00000002",
  1570 => x"00001d44",
  1571 => x"00001155",
  1572 => x"00000002",
  1573 => x"00001d62",
  1574 => x"00001155",
  1575 => x"00000002",
  1576 => x"00001d80",
  1577 => x"00001155",
  1578 => x"00000002",
  1579 => x"00001d9e",
  1580 => x"00001155",
  1581 => x"00000002",
  1582 => x"00001dbc",
  1583 => x"00001155",
  1584 => x"00000002",
  1585 => x"00001dda",
  1586 => x"00001155",
  1587 => x"00000002",
  1588 => x"00001df8",
  1589 => x"00001155",
  1590 => x"00000004",
  1591 => x"00001674",
  1592 => x"00000000",
  1593 => x"00000000",
  1594 => x"00000000",
  1595 => x"000012e7",
  1596 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

