-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbc",
     9 => x"b0080b0b",
    10 => x"0bbcb408",
    11 => x"0b0b0bbc",
    12 => x"b8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bcb80c0b",
    16 => x"0b0bbcb4",
    17 => x"0c0b0b0b",
    18 => x"bcb00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb0e8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bcb07080",
    57 => x"c6e0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e304",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbcc00c",
    65 => x"9f0bbcc4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bcc408ff",
    69 => x"05bcc40c",
    70 => x"bcc40880",
    71 => x"25eb38bc",
    72 => x"c008ff05",
    73 => x"bcc00cbc",
    74 => x"c0088025",
    75 => x"d738800b",
    76 => x"bcc40c80",
    77 => x"0bbcc00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbcc008",
    97 => x"258f3882",
    98 => x"bd2dbcc0",
    99 => x"08ff05bc",
   100 => x"c00c82ff",
   101 => x"04bcc008",
   102 => x"bcc40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bcc008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bcc4",
   111 => x"088105bc",
   112 => x"c40cbcc4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbcc40c",
   116 => x"bcc00881",
   117 => x"05bcc00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bc",
   122 => x"c4088105",
   123 => x"bcc40cbc",
   124 => x"c408a02e",
   125 => x"0981068e",
   126 => x"38800bbc",
   127 => x"c40cbcc0",
   128 => x"088105bc",
   129 => x"c00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbcc8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbcc80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bc",
   169 => x"c8088407",
   170 => x"bcc80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb7b8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bcc80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bcb00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402d0",
   222 => x"050d7d54",
   223 => x"805ba40b",
   224 => x"ec0c7352",
   225 => x"bccc51a8",
   226 => x"892dbcb0",
   227 => x"087b2e81",
   228 => x"ab38bcd0",
   229 => x"0870f80c",
   230 => x"891580f5",
   231 => x"2d8a1680",
   232 => x"f52d7182",
   233 => x"80290588",
   234 => x"1780f52d",
   235 => x"70848080",
   236 => x"2912f40c",
   237 => x"7eff155c",
   238 => x"5e575556",
   239 => x"58767b2e",
   240 => x"8b38811a",
   241 => x"77812a58",
   242 => x"5a76f738",
   243 => x"f71a5a81",
   244 => x"5b807825",
   245 => x"80e63879",
   246 => x"52765184",
   247 => x"8b2dbd98",
   248 => x"52bccc51",
   249 => x"aac82dbc",
   250 => x"b008802e",
   251 => x"b838bd98",
   252 => x"5c83fc59",
   253 => x"7b708405",
   254 => x"5d087081",
   255 => x"ff067188",
   256 => x"2a7081ff",
   257 => x"0673902a",
   258 => x"7081ff06",
   259 => x"75982ae8",
   260 => x"0ce80c58",
   261 => x"e80c57e8",
   262 => x"0cfc1a5a",
   263 => x"53788025",
   264 => x"d33888ac",
   265 => x"04bcb008",
   266 => x"5b848058",
   267 => x"bccc51aa",
   268 => x"9a2dfc80",
   269 => x"18811858",
   270 => x"5887d104",
   271 => x"86b72d84",
   272 => x"0bec0c7a",
   273 => x"802e8d38",
   274 => x"b7bc5190",
   275 => x"af2d8eb2",
   276 => x"2d88da04",
   277 => x"ba805190",
   278 => x"af2d7abc",
   279 => x"b00c02b0",
   280 => x"050d0402",
   281 => x"ec050d84",
   282 => x"0bec0c8e",
   283 => x"932d8afd",
   284 => x"2d81f82d",
   285 => x"9efe2dbc",
   286 => x"b008802e",
   287 => x"81ea3886",
   288 => x"f651b0e2",
   289 => x"2db7bc51",
   290 => x"90af2d8e",
   291 => x"b22d8b89",
   292 => x"2d90bf2d",
   293 => x"b7d00b80",
   294 => x"f52d7086",
   295 => x"2b80c006",
   296 => x"b7dc0b80",
   297 => x"f52d7087",
   298 => x"2b818006",
   299 => x"b7e80b80",
   300 => x"f52d7085",
   301 => x"2ba00674",
   302 => x"730707b7",
   303 => x"f40b80f5",
   304 => x"2d708c2b",
   305 => x"80e08006",
   306 => x"b8800b80",
   307 => x"f52d7084",
   308 => x"2b900674",
   309 => x"730707b8",
   310 => x"8c0b80f5",
   311 => x"2d70912b",
   312 => x"98808006",
   313 => x"b8980b80",
   314 => x"f52d708a",
   315 => x"2b988006",
   316 => x"74730707",
   317 => x"b8a40b80",
   318 => x"f52d7090",
   319 => x"2b848080",
   320 => x"06b8b00b",
   321 => x"80f52d70",
   322 => x"8e2b8380",
   323 => x"80067473",
   324 => x"0707b8bc",
   325 => x"0b80f52d",
   326 => x"70932ba0",
   327 => x"808006b8",
   328 => x"c80b80f5",
   329 => x"2d70942b",
   330 => x"90800a06",
   331 => x"74730707",
   332 => x"b8d40b80",
   333 => x"f52d7088",
   334 => x"2b868006",
   335 => x"7207fc0c",
   336 => x"53545454",
   337 => x"54545454",
   338 => x"54545454",
   339 => x"54545454",
   340 => x"56545257",
   341 => x"57535386",
   342 => x"52bcb008",
   343 => x"8538bcb0",
   344 => x"085271ec",
   345 => x"0c898e04",
   346 => x"800bbcb0",
   347 => x"0c029405",
   348 => x"0d047198",
   349 => x"0c04ffb0",
   350 => x"08bcb00c",
   351 => x"04810bff",
   352 => x"b00c0480",
   353 => x"0bffb00c",
   354 => x"0402f405",
   355 => x"0d8c8b04",
   356 => x"bcb00881",
   357 => x"f02e0981",
   358 => x"06893881",
   359 => x"0bbae40c",
   360 => x"8c8b04bc",
   361 => x"b00881e0",
   362 => x"2e098106",
   363 => x"8938810b",
   364 => x"bae80c8c",
   365 => x"8b04bcb0",
   366 => x"0852bae8",
   367 => x"08802e88",
   368 => x"38bcb008",
   369 => x"81800552",
   370 => x"71842c72",
   371 => x"8f065353",
   372 => x"bae40880",
   373 => x"2e993872",
   374 => x"8429baa4",
   375 => x"05721381",
   376 => x"712b7009",
   377 => x"73080673",
   378 => x"0c515353",
   379 => x"8c810472",
   380 => x"8429baa4",
   381 => x"05721383",
   382 => x"712b7208",
   383 => x"07720c53",
   384 => x"53800bba",
   385 => x"e80c800b",
   386 => x"bae40cbc",
   387 => x"d8518d8c",
   388 => x"2dbcb008",
   389 => x"ff24fef8",
   390 => x"38800bbc",
   391 => x"b00c028c",
   392 => x"050d0402",
   393 => x"f8050dba",
   394 => x"a4528f51",
   395 => x"80727084",
   396 => x"05540cff",
   397 => x"11517080",
   398 => x"25f23802",
   399 => x"88050d04",
   400 => x"02f0050d",
   401 => x"75518b83",
   402 => x"2d70822c",
   403 => x"fc06baa4",
   404 => x"1172109e",
   405 => x"06710870",
   406 => x"722a7083",
   407 => x"0682742b",
   408 => x"70097406",
   409 => x"760c5451",
   410 => x"56575351",
   411 => x"538afd2d",
   412 => x"71bcb00c",
   413 => x"0290050d",
   414 => x"0402fc05",
   415 => x"0d725180",
   416 => x"710c800b",
   417 => x"84120c02",
   418 => x"84050d04",
   419 => x"02f0050d",
   420 => x"75700884",
   421 => x"12085353",
   422 => x"53ff5471",
   423 => x"712ea838",
   424 => x"8b832d84",
   425 => x"13087084",
   426 => x"29148811",
   427 => x"70087081",
   428 => x"ff068418",
   429 => x"08811187",
   430 => x"06841a0c",
   431 => x"53515551",
   432 => x"51518afd",
   433 => x"2d715473",
   434 => x"bcb00c02",
   435 => x"90050d04",
   436 => x"02f8050d",
   437 => x"8b832de0",
   438 => x"08708b2a",
   439 => x"70810651",
   440 => x"52527080",
   441 => x"2e9d38bc",
   442 => x"d8087084",
   443 => x"29bce005",
   444 => x"7381ff06",
   445 => x"710c5151",
   446 => x"bcd80881",
   447 => x"118706bc",
   448 => x"d80c5180",
   449 => x"0bbd800c",
   450 => x"8af62d8a",
   451 => x"fd2d0288",
   452 => x"050d0402",
   453 => x"fc050dbc",
   454 => x"d8518cf9",
   455 => x"2d8ca32d",
   456 => x"8dd0518a",
   457 => x"f22d0284",
   458 => x"050d04bd",
   459 => x"8408bcb0",
   460 => x"0c0402fc",
   461 => x"050d8ebc",
   462 => x"048b892d",
   463 => x"80f6518c",
   464 => x"c02dbcb0",
   465 => x"08f33880",
   466 => x"da518cc0",
   467 => x"2dbcb008",
   468 => x"e838bcb0",
   469 => x"08baf00c",
   470 => x"bcb00851",
   471 => x"84f02d02",
   472 => x"84050d04",
   473 => x"02ec050d",
   474 => x"76548052",
   475 => x"870b8815",
   476 => x"80f52d56",
   477 => x"53747224",
   478 => x"8338a053",
   479 => x"725182f9",
   480 => x"2d81128b",
   481 => x"1580f52d",
   482 => x"54527272",
   483 => x"25de3802",
   484 => x"94050d04",
   485 => x"02f0050d",
   486 => x"bd840854",
   487 => x"81f82d80",
   488 => x"0bbd880c",
   489 => x"7308802e",
   490 => x"81803882",
   491 => x"0bbcc40c",
   492 => x"bd88088f",
   493 => x"06bcc00c",
   494 => x"73085271",
   495 => x"832e9638",
   496 => x"71832689",
   497 => x"3871812e",
   498 => x"af389095",
   499 => x"0471852e",
   500 => x"9f389095",
   501 => x"04881480",
   502 => x"f52d8415",
   503 => x"08b68453",
   504 => x"545285fe",
   505 => x"2d718429",
   506 => x"13700852",
   507 => x"52909904",
   508 => x"73518ee4",
   509 => x"2d909504",
   510 => x"baec0888",
   511 => x"15082c70",
   512 => x"81065152",
   513 => x"71802e87",
   514 => x"38b68851",
   515 => x"909204b6",
   516 => x"8c5185fe",
   517 => x"2d841408",
   518 => x"5185fe2d",
   519 => x"bd880881",
   520 => x"05bd880c",
   521 => x"8c14548f",
   522 => x"a4040290",
   523 => x"050d0471",
   524 => x"bd840c8f",
   525 => x"942dbd88",
   526 => x"08ff05bd",
   527 => x"8c0c0402",
   528 => x"e8050dbd",
   529 => x"8408bd90",
   530 => x"08575587",
   531 => x"518cc02d",
   532 => x"bcb00881",
   533 => x"2a708106",
   534 => x"51527180",
   535 => x"2ea03890",
   536 => x"e5048b89",
   537 => x"2d87518c",
   538 => x"c02dbcb0",
   539 => x"08f438ba",
   540 => x"f0088132",
   541 => x"70baf00c",
   542 => x"70525284",
   543 => x"f02d80fe",
   544 => x"518cc02d",
   545 => x"bcb00880",
   546 => x"2ea638ba",
   547 => x"f008802e",
   548 => x"9138800b",
   549 => x"baf00c80",
   550 => x"5184f02d",
   551 => x"91a2048b",
   552 => x"892d80fe",
   553 => x"518cc02d",
   554 => x"bcb008f3",
   555 => x"3886e22d",
   556 => x"baf00890",
   557 => x"3881fd51",
   558 => x"8cc02d81",
   559 => x"fa518cc0",
   560 => x"2d96f504",
   561 => x"81f5518c",
   562 => x"c02dbcb0",
   563 => x"08812a70",
   564 => x"81065152",
   565 => x"71802eaf",
   566 => x"38bd8c08",
   567 => x"5271802e",
   568 => x"8938ff12",
   569 => x"bd8c0c92",
   570 => x"8704bd88",
   571 => x"0810bd88",
   572 => x"08057084",
   573 => x"29165152",
   574 => x"88120880",
   575 => x"2e8938ff",
   576 => x"51881208",
   577 => x"52712d81",
   578 => x"f2518cc0",
   579 => x"2dbcb008",
   580 => x"812a7081",
   581 => x"06515271",
   582 => x"802eb138",
   583 => x"bd8808ff",
   584 => x"11bd8c08",
   585 => x"56535373",
   586 => x"72258938",
   587 => x"8114bd8c",
   588 => x"0c92cc04",
   589 => x"72101370",
   590 => x"84291651",
   591 => x"52881208",
   592 => x"802e8938",
   593 => x"fe518812",
   594 => x"0852712d",
   595 => x"81fd518c",
   596 => x"c02dbcb0",
   597 => x"08812a70",
   598 => x"81065152",
   599 => x"71802ead",
   600 => x"38bd8c08",
   601 => x"802e8938",
   602 => x"800bbd8c",
   603 => x"0c938d04",
   604 => x"bd880810",
   605 => x"bd880805",
   606 => x"70842916",
   607 => x"51528812",
   608 => x"08802e89",
   609 => x"38fd5188",
   610 => x"12085271",
   611 => x"2d81fa51",
   612 => x"8cc02dbc",
   613 => x"b008812a",
   614 => x"70810651",
   615 => x"5271802e",
   616 => x"ae38bd88",
   617 => x"08ff1154",
   618 => x"52bd8c08",
   619 => x"73258838",
   620 => x"72bd8c0c",
   621 => x"93cf0471",
   622 => x"10127084",
   623 => x"29165152",
   624 => x"88120880",
   625 => x"2e8938fc",
   626 => x"51881208",
   627 => x"52712dbd",
   628 => x"8c087053",
   629 => x"5473802e",
   630 => x"8a388c15",
   631 => x"ff155555",
   632 => x"93d50482",
   633 => x"0bbcc40c",
   634 => x"718f06bc",
   635 => x"c00c81eb",
   636 => x"518cc02d",
   637 => x"bcb00881",
   638 => x"2a708106",
   639 => x"51527180",
   640 => x"2ead3874",
   641 => x"08852e09",
   642 => x"8106a438",
   643 => x"881580f5",
   644 => x"2dff0552",
   645 => x"71881681",
   646 => x"b72d7198",
   647 => x"2b527180",
   648 => x"25883880",
   649 => x"0b881681",
   650 => x"b72d7451",
   651 => x"8ee42d81",
   652 => x"f4518cc0",
   653 => x"2dbcb008",
   654 => x"812a7081",
   655 => x"06515271",
   656 => x"802eb338",
   657 => x"7408852e",
   658 => x"098106aa",
   659 => x"38881580",
   660 => x"f52d8105",
   661 => x"52718816",
   662 => x"81b72d71",
   663 => x"81ff068b",
   664 => x"1680f52d",
   665 => x"54527272",
   666 => x"27873872",
   667 => x"881681b7",
   668 => x"2d74518e",
   669 => x"e42d80da",
   670 => x"518cc02d",
   671 => x"bcb00881",
   672 => x"2a708106",
   673 => x"51527180",
   674 => x"2e81a638",
   675 => x"bd8408bd",
   676 => x"8c085553",
   677 => x"73802e8a",
   678 => x"388c13ff",
   679 => x"15555395",
   680 => x"94047208",
   681 => x"5271822e",
   682 => x"a6387182",
   683 => x"26893871",
   684 => x"812ea938",
   685 => x"96b10471",
   686 => x"832eb138",
   687 => x"71842e09",
   688 => x"810680ed",
   689 => x"38881308",
   690 => x"5190af2d",
   691 => x"96b104bd",
   692 => x"8c085188",
   693 => x"13085271",
   694 => x"2d96b104",
   695 => x"810b8814",
   696 => x"082bbaec",
   697 => x"0832baec",
   698 => x"0c968704",
   699 => x"881380f5",
   700 => x"2d81058b",
   701 => x"1480f52d",
   702 => x"53547174",
   703 => x"24833880",
   704 => x"54738814",
   705 => x"81b72d8f",
   706 => x"942d96b1",
   707 => x"04750880",
   708 => x"2ea23875",
   709 => x"08518cc0",
   710 => x"2dbcb008",
   711 => x"81065271",
   712 => x"802e8b38",
   713 => x"bd8c0851",
   714 => x"84160852",
   715 => x"712d8816",
   716 => x"5675da38",
   717 => x"8054800b",
   718 => x"bcc40c73",
   719 => x"8f06bcc0",
   720 => x"0ca05273",
   721 => x"bd8c082e",
   722 => x"09810698",
   723 => x"38bd8808",
   724 => x"ff057432",
   725 => x"70098105",
   726 => x"7072079f",
   727 => x"2a917131",
   728 => x"51515353",
   729 => x"715182f9",
   730 => x"2d811454",
   731 => x"8e7425c6",
   732 => x"38baf008",
   733 => x"5271bcb0",
   734 => x"0c029805",
   735 => x"0d0402f4",
   736 => x"050dd452",
   737 => x"81ff720c",
   738 => x"71085381",
   739 => x"ff720c72",
   740 => x"882b83fe",
   741 => x"80067208",
   742 => x"7081ff06",
   743 => x"51525381",
   744 => x"ff720c72",
   745 => x"7107882b",
   746 => x"72087081",
   747 => x"ff065152",
   748 => x"5381ff72",
   749 => x"0c727107",
   750 => x"882b7208",
   751 => x"7081ff06",
   752 => x"7207bcb0",
   753 => x"0c525302",
   754 => x"8c050d04",
   755 => x"02f4050d",
   756 => x"74767181",
   757 => x"ff06d40c",
   758 => x"5353bd94",
   759 => x"08853871",
   760 => x"892b5271",
   761 => x"982ad40c",
   762 => x"71902a70",
   763 => x"81ff06d4",
   764 => x"0c517188",
   765 => x"2a7081ff",
   766 => x"06d40c51",
   767 => x"7181ff06",
   768 => x"d40c7290",
   769 => x"2a7081ff",
   770 => x"06d40c51",
   771 => x"d4087081",
   772 => x"ff065151",
   773 => x"82b8bf52",
   774 => x"7081ff2e",
   775 => x"09810694",
   776 => x"3881ff0b",
   777 => x"d40cd408",
   778 => x"7081ff06",
   779 => x"ff145451",
   780 => x"5171e538",
   781 => x"70bcb00c",
   782 => x"028c050d",
   783 => x"0402fc05",
   784 => x"0d81c751",
   785 => x"81ff0bd4",
   786 => x"0cff1151",
   787 => x"708025f4",
   788 => x"38028405",
   789 => x"0d0402f4",
   790 => x"050d81ff",
   791 => x"0bd40c93",
   792 => x"53805287",
   793 => x"fc80c151",
   794 => x"97cc2dbc",
   795 => x"b0088b38",
   796 => x"81ff0bd4",
   797 => x"0c815399",
   798 => x"830498bd",
   799 => x"2dff1353",
   800 => x"72df3872",
   801 => x"bcb00c02",
   802 => x"8c050d04",
   803 => x"02ec050d",
   804 => x"810bbd94",
   805 => x"0c8454d0",
   806 => x"08708f2a",
   807 => x"70810651",
   808 => x"515372f3",
   809 => x"3872d00c",
   810 => x"98bd2db6",
   811 => x"905185fe",
   812 => x"2dd00870",
   813 => x"8f2a7081",
   814 => x"06515153",
   815 => x"72f33881",
   816 => x"0bd00cb1",
   817 => x"53805284",
   818 => x"d480c051",
   819 => x"97cc2dbc",
   820 => x"b008812e",
   821 => x"93387282",
   822 => x"2ebd38ff",
   823 => x"135372e5",
   824 => x"38ff1454",
   825 => x"73ffb038",
   826 => x"98bd2d83",
   827 => x"aa52849c",
   828 => x"80c85197",
   829 => x"cc2dbcb0",
   830 => x"08812e09",
   831 => x"81069238",
   832 => x"96fe2dbc",
   833 => x"b00883ff",
   834 => x"ff065372",
   835 => x"83aa2e9d",
   836 => x"3898d62d",
   837 => x"9aa804b6",
   838 => x"9c5185fe",
   839 => x"2d80539b",
   840 => x"f604b6b4",
   841 => x"5185fe2d",
   842 => x"80549bc8",
   843 => x"0481ff0b",
   844 => x"d40cb154",
   845 => x"98bd2d8f",
   846 => x"cf538052",
   847 => x"87fc80f7",
   848 => x"5197cc2d",
   849 => x"bcb00855",
   850 => x"bcb00881",
   851 => x"2e098106",
   852 => x"9b3881ff",
   853 => x"0bd40c82",
   854 => x"0a52849c",
   855 => x"80e95197",
   856 => x"cc2dbcb0",
   857 => x"08802e8d",
   858 => x"3898bd2d",
   859 => x"ff135372",
   860 => x"c9389bbb",
   861 => x"0481ff0b",
   862 => x"d40cbcb0",
   863 => x"085287fc",
   864 => x"80fa5197",
   865 => x"cc2dbcb0",
   866 => x"08b13881",
   867 => x"ff0bd40c",
   868 => x"d4085381",
   869 => x"ff0bd40c",
   870 => x"81ff0bd4",
   871 => x"0c81ff0b",
   872 => x"d40c81ff",
   873 => x"0bd40c72",
   874 => x"862a7081",
   875 => x"06765651",
   876 => x"53729538",
   877 => x"bcb00854",
   878 => x"9bc80473",
   879 => x"822efee2",
   880 => x"38ff1454",
   881 => x"73feed38",
   882 => x"73bd940c",
   883 => x"738b3881",
   884 => x"5287fc80",
   885 => x"d05197cc",
   886 => x"2d81ff0b",
   887 => x"d40cd008",
   888 => x"708f2a70",
   889 => x"81065151",
   890 => x"5372f338",
   891 => x"72d00c81",
   892 => x"ff0bd40c",
   893 => x"815372bc",
   894 => x"b00c0294",
   895 => x"050d0402",
   896 => x"e8050d78",
   897 => x"55805681",
   898 => x"ff0bd40c",
   899 => x"d008708f",
   900 => x"2a708106",
   901 => x"51515372",
   902 => x"f3388281",
   903 => x"0bd00c81",
   904 => x"ff0bd40c",
   905 => x"775287fc",
   906 => x"80d15197",
   907 => x"cc2d80db",
   908 => x"c6df54bc",
   909 => x"b008802e",
   910 => x"8a38b6d4",
   911 => x"5185fe2d",
   912 => x"9d960481",
   913 => x"ff0bd40c",
   914 => x"d4087081",
   915 => x"ff065153",
   916 => x"7281fe2e",
   917 => x"0981069d",
   918 => x"3880ff53",
   919 => x"96fe2dbc",
   920 => x"b0087570",
   921 => x"8405570c",
   922 => x"ff135372",
   923 => x"8025ed38",
   924 => x"81569cfb",
   925 => x"04ff1454",
   926 => x"73c93881",
   927 => x"ff0bd40c",
   928 => x"81ff0bd4",
   929 => x"0cd00870",
   930 => x"8f2a7081",
   931 => x"06515153",
   932 => x"72f33872",
   933 => x"d00c75bc",
   934 => x"b00c0298",
   935 => x"050d0402",
   936 => x"e8050d77",
   937 => x"797b5855",
   938 => x"55805372",
   939 => x"7625a338",
   940 => x"74708105",
   941 => x"5680f52d",
   942 => x"74708105",
   943 => x"5680f52d",
   944 => x"52527171",
   945 => x"2e863881",
   946 => x"519dd404",
   947 => x"8113539d",
   948 => x"ab048051",
   949 => x"70bcb00c",
   950 => x"0298050d",
   951 => x"0402ec05",
   952 => x"0d765574",
   953 => x"802ebe38",
   954 => x"9a1580e0",
   955 => x"2d51aba1",
   956 => x"2dbcb008",
   957 => x"bcb00880",
   958 => x"c3c80cbc",
   959 => x"b0085454",
   960 => x"80c3a408",
   961 => x"802e9938",
   962 => x"941580e0",
   963 => x"2d51aba1",
   964 => x"2dbcb008",
   965 => x"902b83ff",
   966 => x"f00a0670",
   967 => x"75075153",
   968 => x"7280c3c8",
   969 => x"0c80c3c8",
   970 => x"08537280",
   971 => x"2e9d3880",
   972 => x"c39c08fe",
   973 => x"14712980",
   974 => x"c3b00805",
   975 => x"80c3cc0c",
   976 => x"70842b80",
   977 => x"c3a80c54",
   978 => x"9ef90480",
   979 => x"c3b40880",
   980 => x"c3c80c80",
   981 => x"c3b80880",
   982 => x"c3cc0c80",
   983 => x"c3a40880",
   984 => x"2e8b3880",
   985 => x"c39c0884",
   986 => x"2b539ef4",
   987 => x"0480c3bc",
   988 => x"08842b53",
   989 => x"7280c3a8",
   990 => x"0c029405",
   991 => x"0d0402d8",
   992 => x"050d800b",
   993 => x"80c3a40c",
   994 => x"8454998c",
   995 => x"2dbcb008",
   996 => x"802e9538",
   997 => x"bd985280",
   998 => x"519bff2d",
   999 => x"bcb00880",
  1000 => x"2e8638fe",
  1001 => x"549fb004",
  1002 => x"ff145473",
  1003 => x"8024db38",
  1004 => x"738c38b6",
  1005 => x"e45185fe",
  1006 => x"2d7355a4",
  1007 => x"da048056",
  1008 => x"810b80c3",
  1009 => x"d00c8853",
  1010 => x"b6f852bd",
  1011 => x"ce519d9f",
  1012 => x"2dbcb008",
  1013 => x"762e0981",
  1014 => x"068838bc",
  1015 => x"b00880c3",
  1016 => x"d00c8853",
  1017 => x"b78452bd",
  1018 => x"ea519d9f",
  1019 => x"2dbcb008",
  1020 => x"8838bcb0",
  1021 => x"0880c3d0",
  1022 => x"0c80c3d0",
  1023 => x"08802e80",
  1024 => x"fc3880c0",
  1025 => x"de0b80f5",
  1026 => x"2d80c0df",
  1027 => x"0b80f52d",
  1028 => x"71982b71",
  1029 => x"902b0780",
  1030 => x"c0e00b80",
  1031 => x"f52d7088",
  1032 => x"2b720780",
  1033 => x"c0e10b80",
  1034 => x"f52d7107",
  1035 => x"80c1960b",
  1036 => x"80f52d80",
  1037 => x"c1970b80",
  1038 => x"f52d7188",
  1039 => x"2b07535f",
  1040 => x"54525a56",
  1041 => x"57557381",
  1042 => x"abaa2e09",
  1043 => x"81068d38",
  1044 => x"7551aaf1",
  1045 => x"2dbcb008",
  1046 => x"56a0e904",
  1047 => x"7382d4d5",
  1048 => x"2e8738b7",
  1049 => x"9051a1ab",
  1050 => x"04bd9852",
  1051 => x"75519bff",
  1052 => x"2dbcb008",
  1053 => x"55bcb008",
  1054 => x"802e83de",
  1055 => x"388853b7",
  1056 => x"8452bdea",
  1057 => x"519d9f2d",
  1058 => x"bcb0088a",
  1059 => x"38810b80",
  1060 => x"c3a40ca1",
  1061 => x"b1048853",
  1062 => x"b6f852bd",
  1063 => x"ce519d9f",
  1064 => x"2dbcb008",
  1065 => x"802e8a38",
  1066 => x"b7a45185",
  1067 => x"fe2da28d",
  1068 => x"0480c196",
  1069 => x"0b80f52d",
  1070 => x"547380d5",
  1071 => x"2e098106",
  1072 => x"80cb3880",
  1073 => x"c1970b80",
  1074 => x"f52d5473",
  1075 => x"81aa2e09",
  1076 => x"8106ba38",
  1077 => x"800bbd98",
  1078 => x"0b80f52d",
  1079 => x"56547481",
  1080 => x"e92e8338",
  1081 => x"81547481",
  1082 => x"eb2e8c38",
  1083 => x"80557375",
  1084 => x"2e098106",
  1085 => x"82e438bd",
  1086 => x"a30b80f5",
  1087 => x"2d55748d",
  1088 => x"38bda40b",
  1089 => x"80f52d54",
  1090 => x"73822e86",
  1091 => x"388055a4",
  1092 => x"da04bda5",
  1093 => x"0b80f52d",
  1094 => x"7080c39c",
  1095 => x"0cff0580",
  1096 => x"c3a00cbd",
  1097 => x"a60b80f5",
  1098 => x"2dbda70b",
  1099 => x"80f52d58",
  1100 => x"76057782",
  1101 => x"80290570",
  1102 => x"80c3ac0c",
  1103 => x"bda80b80",
  1104 => x"f52d7080",
  1105 => x"c3c00c80",
  1106 => x"c3a40859",
  1107 => x"57587680",
  1108 => x"2e81ac38",
  1109 => x"8853b784",
  1110 => x"52bdea51",
  1111 => x"9d9f2dbc",
  1112 => x"b00881f6",
  1113 => x"3880c39c",
  1114 => x"0870842b",
  1115 => x"80c3a80c",
  1116 => x"7080c3bc",
  1117 => x"0cbdbd0b",
  1118 => x"80f52dbd",
  1119 => x"bc0b80f5",
  1120 => x"2d718280",
  1121 => x"2905bdbe",
  1122 => x"0b80f52d",
  1123 => x"70848080",
  1124 => x"2912bdbf",
  1125 => x"0b80f52d",
  1126 => x"7081800a",
  1127 => x"29127080",
  1128 => x"c3c40c80",
  1129 => x"c3c00871",
  1130 => x"2980c3ac",
  1131 => x"08057080",
  1132 => x"c3b00cbd",
  1133 => x"c50b80f5",
  1134 => x"2dbdc40b",
  1135 => x"80f52d71",
  1136 => x"82802905",
  1137 => x"bdc60b80",
  1138 => x"f52d7084",
  1139 => x"80802912",
  1140 => x"bdc70b80",
  1141 => x"f52d7098",
  1142 => x"2b81f00a",
  1143 => x"06720570",
  1144 => x"80c3b40c",
  1145 => x"fe117e29",
  1146 => x"770580c3",
  1147 => x"b80c5259",
  1148 => x"5243545e",
  1149 => x"51525952",
  1150 => x"5d575957",
  1151 => x"a4d304bd",
  1152 => x"aa0b80f5",
  1153 => x"2dbda90b",
  1154 => x"80f52d71",
  1155 => x"82802905",
  1156 => x"7080c3a8",
  1157 => x"0c70a029",
  1158 => x"83ff0570",
  1159 => x"892a7080",
  1160 => x"c3bc0cbd",
  1161 => x"af0b80f5",
  1162 => x"2dbdae0b",
  1163 => x"80f52d71",
  1164 => x"82802905",
  1165 => x"7080c3c4",
  1166 => x"0c7b7129",
  1167 => x"1e7080c3",
  1168 => x"b80c7d80",
  1169 => x"c3b40c73",
  1170 => x"0580c3b0",
  1171 => x"0c555e51",
  1172 => x"51555580",
  1173 => x"519ddd2d",
  1174 => x"815574bc",
  1175 => x"b00c02a8",
  1176 => x"050d0402",
  1177 => x"ec050d76",
  1178 => x"70872c71",
  1179 => x"80ff0655",
  1180 => x"565480c3",
  1181 => x"a4088a38",
  1182 => x"73882c74",
  1183 => x"81ff0654",
  1184 => x"55bd9852",
  1185 => x"80c3ac08",
  1186 => x"15519bff",
  1187 => x"2dbcb008",
  1188 => x"54bcb008",
  1189 => x"802eb438",
  1190 => x"80c3a408",
  1191 => x"802e9838",
  1192 => x"728429bd",
  1193 => x"98057008",
  1194 => x"5253aaf1",
  1195 => x"2dbcb008",
  1196 => x"f00a0653",
  1197 => x"a5c90472",
  1198 => x"10bd9805",
  1199 => x"7080e02d",
  1200 => x"5253aba1",
  1201 => x"2dbcb008",
  1202 => x"53725473",
  1203 => x"bcb00c02",
  1204 => x"94050d04",
  1205 => x"02e0050d",
  1206 => x"7970842c",
  1207 => x"80c3cc08",
  1208 => x"05718f06",
  1209 => x"52555372",
  1210 => x"8938bd98",
  1211 => x"5273519b",
  1212 => x"ff2d72a0",
  1213 => x"29bd9805",
  1214 => x"54807480",
  1215 => x"f52d5653",
  1216 => x"74732e83",
  1217 => x"38815374",
  1218 => x"81e52e81",
  1219 => x"f1388170",
  1220 => x"74065458",
  1221 => x"72802e81",
  1222 => x"e5388b14",
  1223 => x"80f52d70",
  1224 => x"832a7906",
  1225 => x"58567699",
  1226 => x"38baf408",
  1227 => x"53728938",
  1228 => x"7280c198",
  1229 => x"0b81b72d",
  1230 => x"76baf40c",
  1231 => x"7353a880",
  1232 => x"04758f2e",
  1233 => x"09810681",
  1234 => x"b538749f",
  1235 => x"068d2980",
  1236 => x"c18b1151",
  1237 => x"53811480",
  1238 => x"f52d7370",
  1239 => x"81055581",
  1240 => x"b72d8314",
  1241 => x"80f52d73",
  1242 => x"70810555",
  1243 => x"81b72d85",
  1244 => x"1480f52d",
  1245 => x"73708105",
  1246 => x"5581b72d",
  1247 => x"871480f5",
  1248 => x"2d737081",
  1249 => x"055581b7",
  1250 => x"2d891480",
  1251 => x"f52d7370",
  1252 => x"81055581",
  1253 => x"b72d8e14",
  1254 => x"80f52d73",
  1255 => x"70810555",
  1256 => x"81b72d90",
  1257 => x"1480f52d",
  1258 => x"73708105",
  1259 => x"5581b72d",
  1260 => x"921480f5",
  1261 => x"2d737081",
  1262 => x"055581b7",
  1263 => x"2d941480",
  1264 => x"f52d7370",
  1265 => x"81055581",
  1266 => x"b72d9614",
  1267 => x"80f52d73",
  1268 => x"70810555",
  1269 => x"81b72d98",
  1270 => x"1480f52d",
  1271 => x"73708105",
  1272 => x"5581b72d",
  1273 => x"9c1480f5",
  1274 => x"2d737081",
  1275 => x"055581b7",
  1276 => x"2d9e1480",
  1277 => x"f52d7381",
  1278 => x"b72d77ba",
  1279 => x"f40c8053",
  1280 => x"72bcb00c",
  1281 => x"02a0050d",
  1282 => x"0402cc05",
  1283 => x"0d7e605e",
  1284 => x"5a800b80",
  1285 => x"c3c80880",
  1286 => x"c3cc0859",
  1287 => x"5c568058",
  1288 => x"80c3a808",
  1289 => x"782e81b0",
  1290 => x"38778f06",
  1291 => x"a0175754",
  1292 => x"738f38bd",
  1293 => x"98527651",
  1294 => x"8117579b",
  1295 => x"ff2dbd98",
  1296 => x"56807680",
  1297 => x"f52d5654",
  1298 => x"74742e83",
  1299 => x"38815474",
  1300 => x"81e52e80",
  1301 => x"f7388170",
  1302 => x"7506555c",
  1303 => x"73802e80",
  1304 => x"eb388b16",
  1305 => x"80f52d98",
  1306 => x"06597880",
  1307 => x"df388b53",
  1308 => x"7c527551",
  1309 => x"9d9f2dbc",
  1310 => x"b00880d0",
  1311 => x"389c1608",
  1312 => x"51aaf12d",
  1313 => x"bcb00884",
  1314 => x"1b0c9a16",
  1315 => x"80e02d51",
  1316 => x"aba12dbc",
  1317 => x"b008bcb0",
  1318 => x"08881c0c",
  1319 => x"bcb00855",
  1320 => x"5580c3a4",
  1321 => x"08802e98",
  1322 => x"38941680",
  1323 => x"e02d51ab",
  1324 => x"a12dbcb0",
  1325 => x"08902b83",
  1326 => x"fff00a06",
  1327 => x"70165154",
  1328 => x"73881b0c",
  1329 => x"787a0c7b",
  1330 => x"54aa9104",
  1331 => x"81185880",
  1332 => x"c3a80878",
  1333 => x"26fed238",
  1334 => x"80c3a408",
  1335 => x"802eb038",
  1336 => x"7a51a4e3",
  1337 => x"2dbcb008",
  1338 => x"bcb00880",
  1339 => x"fffffff8",
  1340 => x"06555b73",
  1341 => x"80ffffff",
  1342 => x"f82e9438",
  1343 => x"bcb008fe",
  1344 => x"0580c39c",
  1345 => x"082980c3",
  1346 => x"b0080557",
  1347 => x"a89e0480",
  1348 => x"5473bcb0",
  1349 => x"0c02b405",
  1350 => x"0d0402f4",
  1351 => x"050d7470",
  1352 => x"08810571",
  1353 => x"0c700880",
  1354 => x"c3a00806",
  1355 => x"5353718e",
  1356 => x"38881308",
  1357 => x"51a4e32d",
  1358 => x"bcb00888",
  1359 => x"140c810b",
  1360 => x"bcb00c02",
  1361 => x"8c050d04",
  1362 => x"02f0050d",
  1363 => x"75881108",
  1364 => x"fe0580c3",
  1365 => x"9c082980",
  1366 => x"c3b00811",
  1367 => x"720880c3",
  1368 => x"a0080605",
  1369 => x"79555354",
  1370 => x"549bff2d",
  1371 => x"0290050d",
  1372 => x"0402f405",
  1373 => x"0d747088",
  1374 => x"2a83fe80",
  1375 => x"06707298",
  1376 => x"2a077288",
  1377 => x"2b87fc80",
  1378 => x"80067398",
  1379 => x"2b81f00a",
  1380 => x"06717307",
  1381 => x"07bcb00c",
  1382 => x"56515351",
  1383 => x"028c050d",
  1384 => x"0402f805",
  1385 => x"0d028e05",
  1386 => x"80f52d74",
  1387 => x"882b0770",
  1388 => x"83ffff06",
  1389 => x"bcb00c51",
  1390 => x"0288050d",
  1391 => x"0402f405",
  1392 => x"0d747678",
  1393 => x"53545280",
  1394 => x"71259738",
  1395 => x"72708105",
  1396 => x"5480f52d",
  1397 => x"72708105",
  1398 => x"5481b72d",
  1399 => x"ff115170",
  1400 => x"eb388072",
  1401 => x"81b72d02",
  1402 => x"8c050d04",
  1403 => x"02e8050d",
  1404 => x"77568070",
  1405 => x"56547376",
  1406 => x"24b33880",
  1407 => x"c3a80874",
  1408 => x"2eab3873",
  1409 => x"51a5d42d",
  1410 => x"bcb008bc",
  1411 => x"b0080981",
  1412 => x"0570bcb0",
  1413 => x"08079f2a",
  1414 => x"77058117",
  1415 => x"57575353",
  1416 => x"74762489",
  1417 => x"3880c3a8",
  1418 => x"087426d7",
  1419 => x"3872bcb0",
  1420 => x"0c029805",
  1421 => x"0d0402f0",
  1422 => x"050dbcac",
  1423 => x"081651ab",
  1424 => x"ec2dbcb0",
  1425 => x"08802e9e",
  1426 => x"388b53bc",
  1427 => x"b0085280",
  1428 => x"c19851ab",
  1429 => x"bd2d80c3",
  1430 => x"d4085473",
  1431 => x"802e8738",
  1432 => x"80c19851",
  1433 => x"732d0290",
  1434 => x"050d0402",
  1435 => x"dc050d80",
  1436 => x"705a5574",
  1437 => x"bcac0825",
  1438 => x"b13880c3",
  1439 => x"a808752e",
  1440 => x"a9387851",
  1441 => x"a5d42dbc",
  1442 => x"b0080981",
  1443 => x"0570bcb0",
  1444 => x"08079f2a",
  1445 => x"7605811b",
  1446 => x"5b565474",
  1447 => x"bcac0825",
  1448 => x"893880c3",
  1449 => x"a8087926",
  1450 => x"d9388055",
  1451 => x"7880c3a8",
  1452 => x"082781d4",
  1453 => x"387851a5",
  1454 => x"d42dbcb0",
  1455 => x"08802e81",
  1456 => x"a838bcb0",
  1457 => x"088b0580",
  1458 => x"f52d7084",
  1459 => x"2a708106",
  1460 => x"77107884",
  1461 => x"2b80c198",
  1462 => x"0b80f52d",
  1463 => x"5c5c5351",
  1464 => x"55567380",
  1465 => x"2e80c938",
  1466 => x"7416822b",
  1467 => x"afac0bbb",
  1468 => x"80120c54",
  1469 => x"77753110",
  1470 => x"80c3d811",
  1471 => x"55569074",
  1472 => x"70810556",
  1473 => x"81b72da0",
  1474 => x"7481b72d",
  1475 => x"7681ff06",
  1476 => x"81165854",
  1477 => x"73802e8a",
  1478 => x"389c5380",
  1479 => x"c19852ae",
  1480 => x"a8048b53",
  1481 => x"bcb00852",
  1482 => x"80c3da16",
  1483 => x"51aee104",
  1484 => x"7416822b",
  1485 => x"acb60bbb",
  1486 => x"80120c54",
  1487 => x"7681ff06",
  1488 => x"81165854",
  1489 => x"73802e8a",
  1490 => x"389c5380",
  1491 => x"c19852ae",
  1492 => x"d8048b53",
  1493 => x"bcb00852",
  1494 => x"77753110",
  1495 => x"80c3d805",
  1496 => x"517655ab",
  1497 => x"bd2daefd",
  1498 => x"04749029",
  1499 => x"75317010",
  1500 => x"80c3d805",
  1501 => x"5154bcb0",
  1502 => x"087481b7",
  1503 => x"2d811959",
  1504 => x"748b24a3",
  1505 => x"38adac04",
  1506 => x"74902975",
  1507 => x"31701080",
  1508 => x"c3d8058c",
  1509 => x"77315751",
  1510 => x"54807481",
  1511 => x"b72d9e14",
  1512 => x"ff165654",
  1513 => x"74f33802",
  1514 => x"a4050d04",
  1515 => x"02fc050d",
  1516 => x"bcac0813",
  1517 => x"51abec2d",
  1518 => x"bcb00880",
  1519 => x"2e8838bc",
  1520 => x"b008519d",
  1521 => x"dd2d800b",
  1522 => x"bcac0cac",
  1523 => x"eb2d8f94",
  1524 => x"2d028405",
  1525 => x"0d0402fc",
  1526 => x"050d7251",
  1527 => x"70fd2ead",
  1528 => x"3870fd24",
  1529 => x"8a3870fc",
  1530 => x"2e80c438",
  1531 => x"b0b70470",
  1532 => x"fe2eb138",
  1533 => x"70ff2e09",
  1534 => x"8106bc38",
  1535 => x"bcac0851",
  1536 => x"70802eb3",
  1537 => x"38ff11bc",
  1538 => x"ac0cb0b7",
  1539 => x"04bcac08",
  1540 => x"f00570bc",
  1541 => x"ac0c5170",
  1542 => x"80259c38",
  1543 => x"800bbcac",
  1544 => x"0cb0b704",
  1545 => x"bcac0881",
  1546 => x"05bcac0c",
  1547 => x"b0b704bc",
  1548 => x"ac089005",
  1549 => x"bcac0cac",
  1550 => x"eb2d8f94",
  1551 => x"2d028405",
  1552 => x"0d0402fc",
  1553 => x"050d800b",
  1554 => x"bcac0cac",
  1555 => x"eb2d8eab",
  1556 => x"2dbcb008",
  1557 => x"bc9c0cba",
  1558 => x"f85190af",
  1559 => x"2d028405",
  1560 => x"0d047180",
  1561 => x"c3d40c04",
  1562 => x"00ffffff",
  1563 => x"ff00ffff",
  1564 => x"ffff00ff",
  1565 => x"ffffff00",
  1566 => x"52657365",
  1567 => x"74000000",
  1568 => x"43617267",
  1569 => x"6172204d",
  1570 => x"6564696f",
  1571 => x"20100000",
  1572 => x"45786974",
  1573 => x"00000000",
  1574 => x"4a6f7973",
  1575 => x"7469636b",
  1576 => x"20437572",
  1577 => x"736f7200",
  1578 => x"4a6f7973",
  1579 => x"7469636b",
  1580 => x"2053696e",
  1581 => x"636c6169",
  1582 => x"72000000",
  1583 => x"4a6f7973",
  1584 => x"7469636b",
  1585 => x"205a5838",
  1586 => x"31000000",
  1587 => x"4368726f",
  1588 => x"6d613831",
  1589 => x"20446573",
  1590 => x"61637469",
  1591 => x"7661646f",
  1592 => x"00000000",
  1593 => x"4368726f",
  1594 => x"6d613831",
  1595 => x"20416374",
  1596 => x"69766164",
  1597 => x"6f000000",
  1598 => x"51532043",
  1599 => x"48525320",
  1600 => x"41637469",
  1601 => x"7661646f",
  1602 => x"28463129",
  1603 => x"00000000",
  1604 => x"51532043",
  1605 => x"48525320",
  1606 => x"44657361",
  1607 => x"63746976",
  1608 => x"61646f00",
  1609 => x"43485224",
  1610 => x"3132382f",
  1611 => x"55444720",
  1612 => x"31323820",
  1613 => x"43686172",
  1614 => x"73000000",
  1615 => x"43485224",
  1616 => x"3132382f",
  1617 => x"55444720",
  1618 => x"36342043",
  1619 => x"68617273",
  1620 => x"00000000",
  1621 => x"43485224",
  1622 => x"3132382f",
  1623 => x"55444720",
  1624 => x"44657361",
  1625 => x"63746976",
  1626 => x"61646f00",
  1627 => x"52414d20",
  1628 => x"42616a61",
  1629 => x"204f6666",
  1630 => x"00000000",
  1631 => x"52414d20",
  1632 => x"42616a61",
  1633 => x"20384b42",
  1634 => x"00000000",
  1635 => x"52414d20",
  1636 => x"5072696e",
  1637 => x"63697061",
  1638 => x"6c203136",
  1639 => x"4b420000",
  1640 => x"52414d20",
  1641 => x"5072696e",
  1642 => x"63697061",
  1643 => x"6c203332",
  1644 => x"4b420000",
  1645 => x"52414d20",
  1646 => x"5072696e",
  1647 => x"63697061",
  1648 => x"6c203438",
  1649 => x"4b420000",
  1650 => x"52414d20",
  1651 => x"5072696e",
  1652 => x"63697061",
  1653 => x"6c20314b",
  1654 => x"42000000",
  1655 => x"56656c6f",
  1656 => x"63696461",
  1657 => x"64204f72",
  1658 => x"6967696e",
  1659 => x"616c0000",
  1660 => x"56656c6f",
  1661 => x"63696461",
  1662 => x"64204e6f",
  1663 => x"57616974",
  1664 => x"00000000",
  1665 => x"56656c6f",
  1666 => x"63696461",
  1667 => x"64207832",
  1668 => x"00000000",
  1669 => x"56656c6f",
  1670 => x"63696461",
  1671 => x"64207838",
  1672 => x"00000000",
  1673 => x"5a583831",
  1674 => x"00000000",
  1675 => x"5a583830",
  1676 => x"00000000",
  1677 => x"5363616e",
  1678 => x"6c696e65",
  1679 => x"73204e6f",
  1680 => x"6e650000",
  1681 => x"5363616e",
  1682 => x"6c696e65",
  1683 => x"73204352",
  1684 => x"54203235",
  1685 => x"25000000",
  1686 => x"5363616e",
  1687 => x"6c696e65",
  1688 => x"73204352",
  1689 => x"54203530",
  1690 => x"25000000",
  1691 => x"5363616e",
  1692 => x"6c696e65",
  1693 => x"73204352",
  1694 => x"54203735",
  1695 => x"25000000",
  1696 => x"426f7264",
  1697 => x"65204e65",
  1698 => x"67726f20",
  1699 => x"4f666600",
  1700 => x"426f7264",
  1701 => x"65204e65",
  1702 => x"67726f20",
  1703 => x"4f6e0000",
  1704 => x"56696465",
  1705 => x"6f20496e",
  1706 => x"7665736f",
  1707 => x"204f6666",
  1708 => x"00000000",
  1709 => x"56696465",
  1710 => x"6f20496e",
  1711 => x"7665736f",
  1712 => x"204f6e00",
  1713 => x"56696465",
  1714 => x"6f204672",
  1715 => x"65712035",
  1716 => x"30487a00",
  1717 => x"56696465",
  1718 => x"6f204672",
  1719 => x"65712036",
  1720 => x"30487a00",
  1721 => x"50656e74",
  1722 => x"61676f6e",
  1723 => x"00000000",
  1724 => x"43617267",
  1725 => x"61204661",
  1726 => x"6c6c6964",
  1727 => x"61000000",
  1728 => x"4f4b0000",
  1729 => x"16200000",
  1730 => x"14200000",
  1731 => x"15200000",
  1732 => x"53442069",
  1733 => x"6e69742e",
  1734 => x"2e2e0a00",
  1735 => x"53442063",
  1736 => x"61726420",
  1737 => x"72657365",
  1738 => x"74206661",
  1739 => x"696c6564",
  1740 => x"210a0000",
  1741 => x"53444843",
  1742 => x"20657272",
  1743 => x"6f72210a",
  1744 => x"00000000",
  1745 => x"57726974",
  1746 => x"65206661",
  1747 => x"696c6564",
  1748 => x"0a000000",
  1749 => x"52656164",
  1750 => x"20666169",
  1751 => x"6c65640a",
  1752 => x"00000000",
  1753 => x"43617264",
  1754 => x"20696e69",
  1755 => x"74206661",
  1756 => x"696c6564",
  1757 => x"0a000000",
  1758 => x"46415431",
  1759 => x"36202020",
  1760 => x"00000000",
  1761 => x"46415433",
  1762 => x"32202020",
  1763 => x"00000000",
  1764 => x"4e6f2070",
  1765 => x"61727469",
  1766 => x"74696f6e",
  1767 => x"20736967",
  1768 => x"0a000000",
  1769 => x"42616420",
  1770 => x"70617274",
  1771 => x"0a000000",
  1772 => x"4261636b",
  1773 => x"00000000",
  1774 => x"00000002",
  1775 => x"00000002",
  1776 => x"00001878",
  1777 => x"0000034e",
  1778 => x"00000003",
  1779 => x"00001cf4",
  1780 => x"00000002",
  1781 => x"00000003",
  1782 => x"00001cec",
  1783 => x"00000002",
  1784 => x"00000003",
  1785 => x"00001ce4",
  1786 => x"00000002",
  1787 => x"00000003",
  1788 => x"00001cd4",
  1789 => x"00000004",
  1790 => x"00000003",
  1791 => x"00001ccc",
  1792 => x"00000002",
  1793 => x"00000003",
  1794 => x"00001cbc",
  1795 => x"00000004",
  1796 => x"00000003",
  1797 => x"00001cac",
  1798 => x"00000004",
  1799 => x"00000003",
  1800 => x"00001ca4",
  1801 => x"00000002",
  1802 => x"00000003",
  1803 => x"00001c98",
  1804 => x"00000003",
  1805 => x"00000003",
  1806 => x"00001c90",
  1807 => x"00000002",
  1808 => x"00000003",
  1809 => x"00001c88",
  1810 => x"00000002",
  1811 => x"00000003",
  1812 => x"00001c7c",
  1813 => x"00000003",
  1814 => x"00000002",
  1815 => x"00001880",
  1816 => x"00001842",
  1817 => x"00000002",
  1818 => x"00001890",
  1819 => x"00000732",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00001898",
  1824 => x"000018a8",
  1825 => x"000018bc",
  1826 => x"000018cc",
  1827 => x"000018e4",
  1828 => x"000018f8",
  1829 => x"00001910",
  1830 => x"00001924",
  1831 => x"0000193c",
  1832 => x"00001954",
  1833 => x"0000196c",
  1834 => x"0000197c",
  1835 => x"0000198c",
  1836 => x"000019a0",
  1837 => x"000019b4",
  1838 => x"000019c8",
  1839 => x"000019dc",
  1840 => x"000019f0",
  1841 => x"00001a04",
  1842 => x"00001a14",
  1843 => x"00001a24",
  1844 => x"00001a2c",
  1845 => x"00001a34",
  1846 => x"00001a44",
  1847 => x"00001a58",
  1848 => x"00001a6c",
  1849 => x"00001a80",
  1850 => x"00001a90",
  1851 => x"00001aa0",
  1852 => x"00001ab4",
  1853 => x"00001ac4",
  1854 => x"00001ad4",
  1855 => x"00001ae4",
  1856 => x"00000004",
  1857 => x"00001af0",
  1858 => x"00001d00",
  1859 => x"00000004",
  1860 => x"00001b00",
  1861 => x"00001bbc",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
  1868 => x"00000000",
  1869 => x"00000000",
  1870 => x"00000000",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"00000000",
  1876 => x"00000000",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000002",
  1887 => x"000021d8",
  1888 => x"00001636",
  1889 => x"00000002",
  1890 => x"000021f6",
  1891 => x"00001636",
  1892 => x"00000002",
  1893 => x"00002214",
  1894 => x"00001636",
  1895 => x"00000002",
  1896 => x"00002232",
  1897 => x"00001636",
  1898 => x"00000002",
  1899 => x"00002250",
  1900 => x"00001636",
  1901 => x"00000002",
  1902 => x"0000226e",
  1903 => x"00001636",
  1904 => x"00000002",
  1905 => x"0000228c",
  1906 => x"00001636",
  1907 => x"00000002",
  1908 => x"000022aa",
  1909 => x"00001636",
  1910 => x"00000002",
  1911 => x"000022c8",
  1912 => x"00001636",
  1913 => x"00000002",
  1914 => x"000022e6",
  1915 => x"00001636",
  1916 => x"00000002",
  1917 => x"00002304",
  1918 => x"00001636",
  1919 => x"00000002",
  1920 => x"00002322",
  1921 => x"00001636",
  1922 => x"00000002",
  1923 => x"00002340",
  1924 => x"00001636",
  1925 => x"00000004",
  1926 => x"00001bb0",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"000017d6",
  1931 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

